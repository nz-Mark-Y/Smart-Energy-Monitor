library verilog;
use verilog.vl_types.all;
entity lab3vhdl_vlg_vec_tst is
end lab3vhdl_vlg_vec_tst;
